module  TLD(
    output         [31:0]   TLD
);

    assign TLD = 32'b0;

endmodule