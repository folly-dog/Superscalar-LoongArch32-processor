module CPUID (
    output       [31:0]  CPUID
);
    
    assign CPUID = 32'b0;

endmodule