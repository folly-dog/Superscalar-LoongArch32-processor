module rename (
    ports
);
    
endmodule